clear && iverilog axi_tb.sv && ./a.out
