
`include "../rtl/axi_slave.sv"
`include "../rtl/axi_master.sv"

`include "../rtl/AXI_UART.sv"

`include "../rtl/UART/UART_SRAM_interface.sv"
`include "../rtl/UART/UART_receive_controller.sv"

`include "../rtl/UART/define_state.h"



module axi_tb;

initial $display("Running axi_tb.sv");

/*

logic clk;
logic reset_n;

logic S_AXIS_TVALID;
logic S_AXIS_TREADY;	

logic [31:0] S_AXIS_TDATA;
logic S_AXIS_TLAST;

logic S_AXIS_TID;
logic S_AXIS_TSTRB;
logic S_AXIS_TKEEP;
logic S_AXIS_TDEST;
logic S_AXIS_TUSER;


axi_slave axi_slave(
	.clk(clk),
	.reset_n(reset_n),

	.S_AXIS_TVALID(S_AXIS_TVALID),
	.S_AXIS_TREADY(S_AXIS_TREADY),	
	
	.S_AXIS_TDATA(S_AXIS_TDATA),
	.S_AXIS_TLAST(S_AXIS_TLAST),
	
	.S_AXIS_TID(S_AXIS_TID),
	.S_AXIS_TSTRB(S_AXIS_TSTRB),
	.S_AXIS_TKEEP(S_AXIS_TKEEP),
	.S_AXIS_TDEST(S_AXIS_TDEST),
	.S_AXIS_TUSER(S_AXIS_TUSER)
);


wire M_AXIS_TVALID;
logic M_AXIS_TREADY;	

wire [31:0] M_AXIS_TDATA;
wire M_AXIS_TLAST;

wire M_AXIS_TID;
wire M_AXIS_TSTRB;
wire M_AXIS_TKEEP;
wire M_AXIS_TDEST;
wire M_AXIS_TUSER;


axi_master axi_master(
	.clk(clk),
	.reset_n(reset_n),

	.M_AXIS_TVALID(M_AXIS_TVALID),
	.M_AXIS_TREADY(M_AXIS_TREADY),	
	
	.M_AXIS_TDATA(M_AXIS_TDATA),
	.M_AXIS_TLAST(M_AXIS_TLAST),
	
	.M_AXIS_TID(M_AXIS_TID),
	.M_AXIS_TSTRB(M_AXIS_TSTRB),
	.M_AXIS_TKEEP(M_AXIS_TKEEP),
	.M_AXIS_TDEST(M_AXIS_TDEST),
	.M_AXIS_TUSER(M_AXIS_TUSER)
);
*/


/*	UART PARAMETERS	*/
parameter C_FAMILY = "virtex6";
parameter C_S_AXI_ACLK_FREQ_HZ = 100_000_000;

parameter C_S_AXI_ADDR_WIDTH = 4;
parameter C_S_AXI_DATA_WIDTH = 32;
parameter C_S_AXI_PROTOCOL = "AXI4LITE";

parameter C_BAUDRATE = 9600;
parameter C_DATA_BITS = 8;
parameter C_USE_PARITY = 0;
parameter C_ODD_PARITY = 0;


/*	UART I/O	*/
logic S_AXI_ACLK;								//P1	-	Clock
logic S_AXI_ARESETN;							//P2	-	Reset (active low)
wire Interrupt;								//P3	-	Interrupt


logic [C_S_AXI_ADDR_WIDTH-1:0] S_AXI_AWADDR;	//P4	-	Write Address
logic S_AXI_AWVALID;							//P5	-	Write Valid
wire S_AXI_AWREADY;							//P6	-	Write Ready


logic [C_S_AXI_DATA_WIDTH-1:0] S_AXI_WDATA;		//P7	-	Write Data
logic [C_S_AXI_DATA_WIDTH/8-1:0] S_AXI_WSTB;	//P8	-	Write Strobes
logic S_AXI_WAVLID;								//P9	-	Write Valid
wire S_AXI_WREADY;								//P10	-	Write Ready


wire [1:0] S_AXI_BRESP;						//P11	-	Write Response (Faults/errors)
wire S_AXI_BVALID;								//P12	-	Write Response Valid
logic S_AXI_BREADY;								//P13	-	Write Response Ready


logic [C_S_AXI_ADDR_WIDTH-1:0] S_AXI_ARADDR;	//P14	-	Read Address
logic S_AXI_ARVALID;							//P15	-	Read Address Valid
wire S_AXI_ARREADY;							//P16	-	Read Address Ready



wire [C_S_AXI_ADDR_WIDTH-1:0] S_AXI_RDATA;		//P17	-	Read Data 
wire [1:0] S_AXI_RRESP;						//P18	-	Read Response (Faults/errors)
wire S_AXI_RVALID;								//P19	-	Read Valid
logic S_AXI_RREADY;								//P20	-	Read Ready

logic RX;										//P21	-	Recieve 
wire TX;										//P22	-	Transmit

//======================================================================//

AXI_UART#(
	.C_FAMILY("virtex6"),
	.C_S_AXI_ACLK_FREQ_HZ(100000000),
	
	.C_S_AXI_ADDR_WIDTH(4),
	.C_S_AXI_DATA_WIDTH(32),
	.C_S_AXI_PROTOCOL("AXI4LITE"),

	.C_BAUDRATE(9600),
	.C_DATA_BITS(8),
	.C_USE_PARITY(0),
	.C_ODD_PARITY(0)
)
AXI_UART (
	.S_AXI_ACLK(S_AXI_ACLK),						//P1	-	Clock
	.S_AXI_ARESETN(S_AXI_ARESETN),					//P2	-	Reset (active low)
	.Interrupt(Interrupt),							//P3	-	Interrupt


	.S_AXI_AWADDR(S_AXI_AWADDR),					//P4	-	Write Address
	.S_AXI_AWVALID(S_AXI_AWVALID),					//P5	-	Write Valid
	.S_AXI_AWREADY(S_AXI_AWREADY),					//P6	-	Write Ready


	.S_AXI_WDATA(S_AXI_WDATA),						//P7	-	Write Data
	.S_AXI_WSTB(S_AXI_WSTB),						//P8	-	Write Strobes
	.S_AXI_WAVLID(S_AXI_WAVLID),					//P9	-	Write Valid
	.S_AXI_WREADY(S_AXI_WREADY),						//P10	-	Write Ready


	.S_AXI_BRESP(S_AXI_BRESP),						//P11	-	Write Response (Faults/errors)
	.S_AXI_BVALID(S_AXI_BVALID),					//P12	-	Write Response Valid
	.S_AXI_BREADY(S_AXI_BREADY),					//P13	-	Write Response Ready


	.S_AXI_ARADDR(S_AXI_ARADDR),					//P14	-	Read Address
	.S_AXI_ARVALID(S_AXI_ARVALID),					//P15	-	Read Address Valid
	.S_AXI_ARREADY(S_AXI_ARREADY),					//P16	-	Read Address Ready


	.S_AXI_RDATA(S_AXI_RDATA),						//P17	-	Read Data 
	.S_AXI_RRESP(S_AXI_RRESP),						//P18	-	Read Response (Faults/errors)
	.S_AXI_RVALID(S_AXI_RVALID),					//P19	-	Read Valid
	.S_AXI_RREADY(S_AXI_RREADY),					//P20	-	Read Ready

	.RX(RX),										//P21	-	Recieve 
	.TX(TX)											//P22	-	Transmit
);




always begin
	S_AXI_ACLK<=0; #5; S_AXI_ACLK<=1;
end







initial begin


end





initial begin
	repeat(10000) @(posedge S_AXI_ACLK);
	$display("Testbench duration exhausted (10,000 clocks) ");
	$finish;
end

endmodule
