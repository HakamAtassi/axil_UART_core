

module top
(

);





endmodule

